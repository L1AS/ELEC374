module shr_op(
  input wire[31:0] A_reg, B_reg,
  output wire[31:0] ror_out
);

endmodule