module rol_op (

);

  

endmodule