module full_adder (
    input a, b, Cin, 
    output sum, Cout
);
wire 

half_adder ha1(.a(a), .b(b), .sum())
endmodule